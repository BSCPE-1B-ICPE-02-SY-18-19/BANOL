CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 120 10
149 75 1534 806
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
338 183 465 292
76546066 0
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 976 37 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9998 0 0
2
5.89884e-315 0
0
2 +V
167 294 256 0 1 3
0 7
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3536 0 0
2
43530.4 0
0
7 Pulser~
4 93 306 0 10 12
0 18 19 8 20 0 0 5 5 1
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4597 0 0
2
43530.4 1
0
9 CC 7-Seg~
183 855 90 0 17 19
10 15 14 13 12 11 10 9 21 2
0 0 1 1 1 1 1 2
0
0 0 21104 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3835 0 0
2
43530.4 2
0
9 2-In AND~
219 685 208 0 3 22
0 16 4 17
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3670 0 0
2
43530.4 3
0
9 2-In AND~
219 523 200 0 3 22
0 6 5 16
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5616 0 0
2
43530.4 4
0
6 74112~
219 757 335 0 7 32
0 7 17 8 17 7 22 3
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
9323 0 0
2
43530.4 5
0
6 74112~
219 610 333 0 7 32
0 7 16 8 16 7 23 4
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
317 0 0
2
43530.4 6
0
6 74112~
219 441 336 0 7 32
0 7 6 8 6 7 24 5
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3108 0 0
2
43530.4 7
0
6 74112~
219 294 336 0 7 32
0 7 7 8 7 7 25 6
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2A
21 -62 42 -54
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
4299 0 0
2
43530.4 8
0
6 74LS48
188 959 315 0 14 29
0 3 4 5 6 26 27 9 10 11
12 13 14 15 28
0
0 0 4832 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9672 0 0
2
43530.4 9
0
37
1 9 2 0 0 8320 0 1 4 0 0 4
976 45
976 51
855 51
855 48
0 1 3 0 0 12416 0 0 11 7 0 5
798 299
798 443
894 443
894 279
927 279
0 2 4 0 0 8320 0 0 11 29 0 5
641 297
641 452
902 452
902 288
927 288
0 3 5 0 0 8320 0 0 11 27 0 5
483 300
483 458
908 458
908 297
927 297
0 4 6 0 0 8320 0 0 11 37 0 5
333 300
333 467
915 467
915 306
927 306
0 1 7 0 0 8192 0 0 2 24 0 4
256 300
256 273
294 273
294 265
7 0 3 0 0 0 0 7 0 0 0 2
781 299
811 299
1 0 7 0 0 0 0 2 0 0 12 2
294 265
294 265
0 0 7 0 0 4096 0 0 0 12 15 2
355 265
355 356
1 1 7 0 0 8192 0 8 7 0 0 4
610 270
610 265
757 265
757 272
1 1 7 0 0 8320 0 9 8 0 0 4
441 273
441 265
610 265
610 270
1 1 7 0 0 0 0 10 9 0 0 4
294 273
294 265
441 265
441 273
5 5 7 0 0 0 0 8 7 0 0 4
610 345
610 356
757 356
757 347
5 5 7 0 0 0 0 9 8 0 0 4
441 348
441 356
610 356
610 345
5 5 7 0 0 0 0 10 9 0 0 4
294 348
294 356
441 356
441 348
3 0 8 0 0 12288 0 3 0 0 34 4
117 297
140 297
140 398
242 398
7 7 9 0 0 12416 0 11 4 0 0 5
991 279
1025 279
1025 174
870 174
870 126
8 6 10 0 0 12416 0 11 4 0 0 5
991 288
1020 288
1020 169
864 169
864 126
9 5 11 0 0 12416 0 11 4 0 0 5
991 297
1015 297
1015 164
858 164
858 126
10 4 12 0 0 12416 0 11 4 0 0 5
991 306
1010 306
1010 159
852 159
852 126
11 3 13 0 0 8320 0 11 4 0 0 5
991 315
1005 315
1005 154
846 154
846 126
12 2 14 0 0 8320 0 11 4 0 0 5
991 324
1000 324
1000 149
840 149
840 126
13 1 15 0 0 8320 0 11 4 0 0 5
991 333
995 333
995 144
834 144
834 126
4 2 7 0 0 0 0 10 10 0 0 4
270 318
256 318
256 300
270 300
2 0 16 0 0 4096 0 8 0 0 26 2
586 297
548 297
0 4 16 0 0 4224 0 0 8 28 0 3
548 200
548 315
586 315
2 7 5 0 0 0 0 6 9 0 0 4
499 209
492 209
492 300
465 300
3 1 16 0 0 0 0 6 5 0 0 4
544 200
548 200
548 199
661 199
2 7 4 0 0 0 0 5 8 0 0 4
661 217
652 217
652 297
634 297
2 0 17 0 0 4096 0 7 0 0 31 2
733 299
712 299
3 4 17 0 0 8320 0 5 7 0 0 4
706 208
712 208
712 317
733 317
3 0 8 0 0 0 0 8 0 0 34 3
580 306
554 306
554 399
3 0 8 0 0 0 0 9 0 0 34 3
411 309
397 309
397 399
3 3 8 0 0 12416 0 10 7 0 0 6
264 309
242 309
242 399
702 399
702 308
727 308
1 0 6 0 0 0 0 6 0 0 36 3
499 191
367 191
367 300
4 0 6 0 0 0 0 9 0 0 37 3
417 318
367 318
367 300
7 2 6 0 0 0 0 10 9 0 0 2
318 300
417 300
2
-27 0 0 0 700 0 0 0 0 3 2 1 66
13 Comic Sans MS
0 0 0 28
27 13 329 113
40 20 315 96
28 BANOL,FELIPE JR. S
BSCpE-1B
-21 0 0 0 400 255 0 0 0 3 2 1 66
12 Segoe Script
0 0 0 35
262 123 780 176
273 131 768 164
35 BINARY 4-BIT SYNCHRONOUS UP COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
